module decoder(a,b,e,y0,y1,y2,y3);
	input a,b,e;
	output y0,y1,y2,y3;
	reg y0,y1,y2,y3;
	
	always @ (a or b or e )
	begin
		
	end
endmodule
